property s109;
    nexttime b[->3];
endproperty