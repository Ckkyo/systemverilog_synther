sequence s24;
    a[->0] ##1 !a[+] ##1 b;
endsequence