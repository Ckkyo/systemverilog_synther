property s102;
    not(a[=1] ##1 b[->2] ##1 a);
endproperty