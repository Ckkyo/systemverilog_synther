property s105;
    (b[->1] ) intersect a;
endproperty