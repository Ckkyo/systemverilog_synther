property s121;
    (c[=3] #-# (a[=3:5] within b[->2]));
endproperty