sequence s14;
    a[=3] ##1 b;
endsequence