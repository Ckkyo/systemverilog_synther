property s116;
    (a[*] |-> (a));
endproperty 