property s104;
    c[*2:3] intersect b[*1:2];
endproperty