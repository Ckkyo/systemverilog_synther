property s115;
    (a ##1 d[*0] ##0 b);
endproperty