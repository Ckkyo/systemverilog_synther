property s115;
    a iff b;
endproperty