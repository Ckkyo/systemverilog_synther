property s128;
    c[=3] until_with !b[->2];
endproperty