sequence s27;
    !a[*0:1] ##1 !a[*0:1] ##1 b;
endsequence