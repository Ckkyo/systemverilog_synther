property s113;
    (c |-> a[*0:1] ##1 b);
endproperty