property s125;
    c[*3] until !b[*2];
endproperty