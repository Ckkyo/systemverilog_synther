sequence s5;
    a ##[*] b;
endsequence
