property s117;
    reject_on(a) b;
endproperty