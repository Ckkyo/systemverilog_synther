property s109;
    (b[->1] and a[=1] );
endproperty