sequence s13;
    a[->1:2];
endsequence