property s103;
    (a[=0:$] ##1 b) or (a[=1] ##1 b[->2] ##1 a);
endproperty