property a2;
    a ##1 b|=> d[*2:4] ##1 e ##1 c;
endproperty 