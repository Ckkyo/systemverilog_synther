property s108;
    b[->1] intersect ( a[=1] ##1 d[*0:$]);
endproperty
