property a5;
    a |=> b[*25] ##1 c;
endproperty 