property axi_r_1;
    arvalid_s0 |-> ##[0:2] arready_s0 ##[1:8] rvalid_s0 ##[0:8] rready_s0;
endproperty 