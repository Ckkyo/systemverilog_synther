sequence s18;
    a[=0:$] ##1 b;
endsequence