property s112;
    (c throughout b[->2]);
endproperty