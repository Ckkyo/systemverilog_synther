property s126;
    c[*3] until(c[*3] and !b[*2]);
endproperty