sequence s17;
    first_match(a ##[2:4] b);
endsequence