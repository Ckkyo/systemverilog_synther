sequence s6;
    a ##[+] b;
endsequence
