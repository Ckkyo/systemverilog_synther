property s100;
    a ##1 a[*] ##1 b;
endproperty