property s106;
    b[->1] intersect a[=1];
endproperty