property s30;
    b[->2];
endproperty