property a1;
    a |=> d[*1:3] ##1 e;
endproperty 