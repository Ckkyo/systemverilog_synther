property s117;
    (c ##0 (a intersect b));
endproperty 