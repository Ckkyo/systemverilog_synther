sequence s3;
    a ##1 b;
endsequence
