sequence s2;
    a ##0 b;
endsequence
