property s129;
    always a;
endproperty