sequence s0;
    a;
endsequence
