sequence s23;
    ##0 ##1 !a[*] ##1 b;
endsequence