property s114;
    not(c[=1]);
endproperty