property a1;
    rib_hold_flag_i[->3] within rst[*10];
endproperty