property s110;
    (a[=3:5] and b[->2]) and c[*1:5];
endproperty