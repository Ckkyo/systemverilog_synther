sequence s9;
    a ##1 ##1 ##1 c;
endsequence

