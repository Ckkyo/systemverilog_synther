sequence s21;
    a[=0:0] ##1 b;
endsequence