property a0;
    ctrl_jump_flag_o[->1] within rst[*1:20];
endproperty 