sequence s12;
    b[->3];
endsequence