sequence s29;
    ##1 a[*];
endsequence
