sequence s1;
    !a;
endsequence
