property s118;
    sync_accept_on(a) b;
endproperty