property s132;
    a iff b;
endproperty