sequence s16;
    !a[->0:$] ##1 b;
endsequence