property a4;
    first_match(a ##[2:4] b);
endproperty 