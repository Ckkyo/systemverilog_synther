sequence s20;
    a[->1] ##1 b[->1];
endsequence