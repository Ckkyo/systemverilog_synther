property s118;
    (c[*] |-> (a ##0 b));
endproperty