property s133;
    (a[=0:$] ##1 b) iff (a[=1] ##1 b[->2] ##1 a);
endproperty