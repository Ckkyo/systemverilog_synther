property a0;
    a ##1 b ##1 c |=> d ##1 e;
endproperty 