sequence s11;
    a[->0] ##1 b;
endsequence