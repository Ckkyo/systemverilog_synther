sequence s8;
    ##1 b;
endsequence
