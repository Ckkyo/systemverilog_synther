sequence s7;
    a[*0] ##1 b;
endsequence
