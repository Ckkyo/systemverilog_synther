property s130;
    a implies b;
endproperty