property a3;
    a |=> b[*0:2] ##1 c;
endproperty 