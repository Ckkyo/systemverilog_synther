property s116;
    accept_on(a) b;
endproperty