property s107;
    (a) intersect b[->1];
endproperty
