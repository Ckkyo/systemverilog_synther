property s111;
    (a[=3:5] within b[->2]);
endproperty