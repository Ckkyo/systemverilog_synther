property s123;
    a within c[*10];
endproperty