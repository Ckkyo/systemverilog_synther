property s101;
    a ##1 b[+];
endproperty