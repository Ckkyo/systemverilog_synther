property s114;
    a implies b;
endproperty