sequence s26;
    !a[*] ##1 !a[*] ##1 b;
endsequence