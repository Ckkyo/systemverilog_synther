sequence s15;
    a[=1:2];
endsequence