property s124;
    c until b;
endproperty