sequence s25;
    ##0 b[->1:3] ##0 ##3 a[*] ##1 ##0 !b[+] ##1 c[*3] ##[+] b[->1:$];
endsequence