property s111;
    eventually[2:30] b[->3];
endproperty