sequence s19;
    a[=1:$] ##1 b;
endsequence