property s122;
    (a #=# (a[=3:5] within b[->2]));
endproperty