sequence s28;
    a[*] ##1 !a;
endsequence