property s119;
    sync_reject_on(a) b;
endproperty