property s120;
    (c[=3] |=> (a[=3:5] within b[->2]));
endproperty