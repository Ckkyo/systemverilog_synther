property s131;
    (a[=0:$] ##1 b) implies (a[=1] ##1 b[->2] ##1 a);
endproperty