sequence s10;
    !a[*] ##1 b;
endsequence
