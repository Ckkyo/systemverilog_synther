sequence s4;
    a ##[1:3] b;
endsequence
