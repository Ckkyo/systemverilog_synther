property axi_r_0;
        arvalid_s0 |-> ##[0:64] arready_s0;
endproperty